library verilog;
use verilog.vl_types.all;
entity mccomp_tb is
end mccomp_tb;
