library verilog;
use verilog.vl_types.all;
entity sccomp_tb is
end sccomp_tb;
